
module altpll (
	altpll_0_c0_clk,
	altpll_0_c1_clk,
	clk_clk,
	reset_reset_n);	

	output		altpll_0_c0_clk;
	output		altpll_0_c1_clk;
	input		clk_clk;
	input		reset_reset_n;
endmodule
